�� sr java.util.ArrayListx����a� I sizexp   w   sr model.Pessoa        L emailt Ljava/lang/String;L nomeq ~ L senhaq ~ xpt gomes@gmail.comt Arthur Gomes Severot 1234sq ~ t joao@gmail.comt João Pedrot #12345asq ~ t juniorarthur@gmail.comt Arthur Juniort 12345sq ~ t nalu@gmail.comt Ana Luísa Hofmannt 1234sq ~ t zinalda@gmai.comt Zinalda Pintot 12345sq ~ t zinaldajr@gmail.comt Zinalda Pinto Juniort 122342sq ~ t joao@gmail.comt João Silvat 1234x