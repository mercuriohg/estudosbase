�� sr java.util.ArrayListx����a� I sizexp   w   sr model.Pessoa        L emailt Ljava/lang/String;L nomeq ~ L senhaq ~ xpt gomes@gmail.comt Arthur Gomes Severot 123456sq ~ t gomesarthur@gmail.comt Arthur Gomes Severot 12345678sq ~ t gomesarthur6@gmail.comt Arthur Gomest 	123456789sq ~ t bh27@gmail.comt Bruno Henriquet $12334x