�� sr java.util.ArrayListx����a� I sizexp   w   sr model.Pessoan��
4� I idL emailt Ljava/lang/String;L nomeq ~ L senhaq ~ L senha2q ~ xp   t admin@gmail.comt adminat 123t 123x