�� sr java.util.ArrayListx����a� I sizexp   w   sr model.Pessoa        L emailt Ljava/lang/String;L nomeq ~ L senhaq ~ L senha2q ~ xpt arthur@gmail.comt Arthurt 12345t 12345sq ~ t um@gmail.comt umt 1234t 1234x